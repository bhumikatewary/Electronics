dudjeenufn
  nssndj
